`ifndef FIFO_DEF_SV
`define FIFO_DEF_SV
  `define DATA_WIDTH 8
  `define DEPTH 16
  `define SIZE $clog2(DEPTH)
  `define DIFF 2
`endif
